`timescale 1ns / 1ns
module control_unit(input[30:0] instr,input zero,output reg memwrite,regwrite,alusrc,output reg[2:0] aluctrl,output reg [1:0]immsrc,resultsrc,output pcsrc);
wire[6:0] op = instr[6:0];
wire funct7=instr[30];
wire[2:0] funct3=instr[14:12];
reg jump;
reg branch;
reg[1:0] alu_op;
assign pcsrc=(zero&branch)|jump;
always@(*)
begin
case (op)
'b0000011:
begin
regwrite=1;
immsrc='b00;
alusrc=1;
memwrite=0;
resultsrc=1;
branch=0;
jump=0;
alu_op='b00;
end
'b0100011:
begin
regwrite=0;
immsrc='b01;
alusrc=1;
memwrite=1;
jump=0;
resultsrc=1;
branch=0;
alu_op='b00;
end
'b0110011:
begin
regwrite=1;
immsrc='b01;
alusrc=0;
memwrite=0;
jump=0;
resultsrc=0;
branch=0;
alu_op='b10;
end
'b1100011:
begin
regwrite=0;
immsrc='b10;
alusrc=0;
jump=0;
memwrite=0;
resultsrc=1;
branch=1;
alu_op='b01;
end
'b0010011:
begin
regwrite=1;
immsrc='b00;
alusrc=1;
jump=0;
memwrite=0;
resultsrc=0;
branch=0;
alu_op='b10;
end
'b1101111:
begin
regwrite=1;
immsrc='b11;
alusrc=0;
jump=1;
memwrite=0;
resultsrc='b10;
branch=0;
alu_op='b01;
end
default:
begin
regwrite=1;
immsrc='b01;
alusrc=1;
memwrite=1;
resultsrc='b10;
branch=0;
alu_op='b00;
jump=0;
end
endcase
end
always@(*)
begin
case(alu_op)
'b00:
aluctrl='b000;
'b01:
aluctrl='b001;
'b10:
begin
case(funct3)
'b000:
begin
if(op[5]==1&&funct7==1)
aluctrl='b001;
else
aluctrl='b000;
end
3'b010:aluctrl='b101;
3'b110:aluctrl='b011;
3'b111:aluctrl='b010;
default:aluctrl=0;
endcase
end
default:aluctrl=0;
endcase
end
endmodule
